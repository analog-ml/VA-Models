* Simple Test

Vd d 0 1.8
Vg g 0 1.2
Vs s 0 0
m1 d g s s nmos 

.op
.end
